
`define DELAY 20 
module lhu_testbench();

wire [31:0] result;

reg [31:0] inputx; 



lhu res(inputx, result[31:0]);

initial begin
inputx = 32'b00000101010101111100010111010101;

#`DELAY;

inputx = 32'b00000101010101010000010101010111;

#`DELAY;
end

initial begin
$monitor("time = %2d, INPUT =%32b, OUTPUT=%32b\n", $time, inputx, result);		
end 

 
endmodule